module Datapath();
wire a;


endmodule